for (i = 0; i < 32; i = i+1)
	mem[i] <= 32'b0;
